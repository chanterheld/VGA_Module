library ieee;
use ieee.std_logic_1164.all;

entity mplex2t1_1 is 
	port(	a	: in 	std_logic;
		b	: in	std_logic;
		sel	: in	std_logic;
		q	: out	std_logic
	);
end entity mplex2t1_1;
