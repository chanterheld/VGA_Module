library ieee;
use ieee.std_logic_1164.all;

entity one_adder_3 is
	port(	a	: in	std_logic_vector(2 downto 0);
		sum	: out	std_logic_vector(2 downto 0)
	);
end entity one_adder_3;
