library ieee;
use ieee.std_logic_1164.all;

entity h_add is
 	port(	a	: in 	std_logic;
 		b	: in 	std_logic;
 		s 	: out 	std_logic;
 		c_out 	: out 	std_logic
	);
end entity h_add;
